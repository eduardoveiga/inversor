Inversor
.include 45nm_HP.pm

*Descricao do circuito

**fontes
 Vin in GND PULSE (0 1 0 20p 20p 200p 260p)

**capacitancia de saida
C1 out 0 5f





Vdd vdd GND 1V
M1 out in vdd vdd   PMOS L=45n W=360n
M2 out in GND GND   NMOS L=45n W=180n

.control
run
plot in out
.endc


*Parametros de Simulação
.tran 1p 1000p

*---- Tempo de propagacao
.measure tran tphl_a trig v(in) val=0.5 rise=1 targ V(out) val=0.5 fall=1
.measure tran tplh_a trig v(in) val=0.5 fall=1 targ V(out) val=0.5 rise=1

*---- Tempo de transicao
.measure tran tfall_a trig v(out) val=0.8 fall=1 targ v(out) val=0.2 fall=1
.measure tran trise_a trig v(out) val=0.2 rise=1 targ v(out) val=0.8 rise=1


.end
